`timescale 1ns / 1ps


module Memory_Control #(parameter DATA_WIDTH = 32,
                        ADDRESS_BUS  = 22,
                        ADDRESS_BITS = 15,
                        ENABLE_BITS  = 7,
                        IFM_SIZE     = 32)
    (
    input clk,
    input [DATA_WIDTH-1:0] riscv_data_bus,
    input [ADDRESS_BUS-1:0] riscv_address_bus,
    input initialization_done, 
    
    output conva1_start,
     
    output [3-1:0] conva1_ifm_enable_write,
    
    output [3-1:0] conva1_wm_enable_write,
    output [3-1:0] convb_wm_enable_write,
    output [3-1:0] conva2_wm_enable_write,
    output [84-1:0] fc1_wm_enable_write,
    output [10-1:0] fc2_wm_enable_write,
    
    output conva1_bm_enable_write,
    output [3-1:0] convb_bm_enable_write,
    output conva2_bm_enable_write,
    output fc1_bm_enable_write,
    output fc2_bm_enable_write,
    
    output [DATA_WIDTH-1:0] riscv_data,
    output [ADDRESS_BITS-1:0] riscv_address
    );
   
    reg [113-1:0] enable_write;
    wire [ENABLE_BITS-1:0] address_enable_bits;
    
    assign riscv_data          = riscv_data_bus;
    assign riscv_address       = riscv_address_bus[ADDRESS_BITS-1:0];
    
    assign address_enable_bits = riscv_address_bus[ADDRESS_BUS-1 : ADDRESS_BUS-ENABLE_BITS];
    
    //-----------------------------------//
    //------------ConvA1-----------------//
    //-----------------------------------//   
   

 assign    conva1_start = initialization_done;
    
 
    always @*
    begin
        case(address_enable_bits)
            //WM ConvA1
            7'd1  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;end
            7'd2  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;end
            7'd3  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;end
                                              
            //WM ConvB1                       
            7'd4  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;end
            7'd5  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;end
            7'd6  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;end
                                              
            //WM ConvA2                       
            7'd7  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;end
            7'd8  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;end
            7'd9  : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;end
                                              
            //WM FC 1                         
            7'd10 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;end
            7'd11 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;end
            7'd12 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;end
            7'd13 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;end
            7'd14 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;end
            7'd15 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;end
            7'd16 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;end
            7'd17 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;end
            7'd18 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;end
            7'd19 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;end
            7'd20 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;end
            7'd21 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;end
            7'd22 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;end
            7'd23 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;end
            7'd24 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;end
            7'd25 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;end 
            7'd26 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;end
            7'd27 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;end
            7'd28 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;end
            7'd29 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;end
            7'd30 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;end
            7'd31 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;end
            7'd32 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;end
            7'd33 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;end
            7'd34 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;end
            7'd35 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;end
            7'd36 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;end
            7'd37 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;end
            7'd38 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;end
            7'd39 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;end
            7'd40 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;end
            7'd41 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;end
            7'd42 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;end
            7'd43 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;end
            7'd44 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;end
            7'd45 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;end
            7'd46 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;end
            7'd47 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;end
            7'd48 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;end
            7'd49 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;end
            7'd50 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;end 
            7'd51 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;end
            7'd52 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;end                    
            7'd53 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;end                
            7'd54 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;end                                             
            7'd55 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;end
            7'd56 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;end
            7'd57 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;end
            7'd58 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;end
            7'd59 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;end
            7'd60 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;end
            7'd61 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;end
            7'd62 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;end
            7'd63 : begin enable_write = 113'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;end
            7'd64 : begin enable_write = 113'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;end
            7'd65 : begin enable_write = 113'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;end
            7'd66 : begin enable_write = 113'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;end
            7'd67 : begin enable_write = 113'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;end
            7'd68 : begin enable_write = 113'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;end
            7'd69 : begin enable_write = 113'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;end
            7'd70 : begin enable_write = 113'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd71 : begin enable_write = 113'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd72 : begin enable_write = 113'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd73 : begin enable_write = 113'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd74 : begin enable_write = 113'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd75 : begin enable_write = 113'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;end            
            7'd76 : begin enable_write = 113'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;end  
            7'd77 : begin enable_write = 113'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd78 : begin enable_write = 113'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd79 : begin enable_write = 113'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd80 : begin enable_write = 113'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd81 : begin enable_write = 113'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd82 : begin enable_write = 113'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd83 : begin enable_write = 113'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd84 : begin enable_write = 113'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd85 : begin enable_write = 113'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd86 : begin enable_write = 113'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd87 : begin enable_write = 113'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd88 : begin enable_write = 113'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd89 : begin enable_write = 113'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd90 : begin enable_write = 113'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd91 : begin enable_write = 113'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd92 : begin enable_write = 113'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd93 : begin enable_write = 113'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
                                             
            //WM FC 2                        
            7'd94 : begin enable_write = 113'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd95 : begin enable_write = 113'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd96 : begin enable_write = 113'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd97 : begin enable_write = 113'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd98 : begin enable_write = 113'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd99 : begin enable_write = 113'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd100: begin enable_write = 113'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd101 : begin enable_write= 113'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd102 : begin enable_write= 113'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd103 : begin enable_write= 113'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
                                             
            //Bias                           
            7'd104 : begin enable_write= 113'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd105 : begin enable_write= 113'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd106 : begin enable_write= 113'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd107 : begin enable_write= 113'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd108 : begin enable_write= 113'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end                               
            7'd109 : begin enable_write= 113'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd110 : begin enable_write= 113'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
          
           //IFM Layer 1
            7'd111 : begin enable_write= 113'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end 
            7'd112 : begin enable_write= 113'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
            7'd113 : begin enable_write= 113'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
                                 
           default : begin enable_write =113'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;end
                                              
        endcase                               
    end                                       
                                              
                                              
                                              
    assign conva1_ifm_enable_write = enable_write[112:110]; 
                                              
    assign conva1_wm_enable_write  = enable_write[2:0];
    assign convb_wm_enable_write   = enable_write[5:3];
    assign conva2_wm_enable_write  = enable_write[8:6];
    assign fc1_wm_enable_write     = enable_write[92:9];
    assign fc2_wm_enable_write     = enable_write[102:93];
    
    assign conva1_bm_enable_write  = enable_write[103];
    assign convb_bm_enable_write   = enable_write[106:104];
    assign conva2_bm_enable_write  = enable_write[107];
    assign fc1_bm_enable_write     = enable_write[108];
    assign fc2_bm_enable_write     = enable_write[109];
    
endmodule
