`timescale 1ns / 1ps


module ConvA2_tb;
    reg clk;
	reg reset;
	reg [31:0] riscv_data_bus;
	reg [17:0] riscv_address_bus;
	reg [31:0] data_in_from_previous;
	reg [7:0] ifm_address_write_previous;
	reg ifm_enable_write_previous;
	reg start_from_previous;
	reg end_from_next;
    reg data_in_from_next;
	// Outputs
	wire end_to_pervious;
	wire [31:0] data_out_for_next;
	//wire [4:0] ifm_address_write_next;
	wire ifm_enable_write_next;
	wire ifm_enable_read_next;
	wire start_to_next;

	// Instantiate the Unit Under Test (UUT)
	TOP_ConvA2 uut (
		.clk(clk), 
		.reset(reset), 
		.riscv_data_bus(riscv_data_bus), 
		.riscv_address_bus(riscv_address_bus), 
		.data_in_from_previous(data_in_from_previous), 
		.ifm_address_write_previous(ifm_address_write_previous), 
		.ifm_enable_write_previous(ifm_enable_write_previous), 
		.start_from_previous(start_from_previous), 
		.end_to_previous(end_to_previous), 
		.end_from_next(end_from_next), 
		.data_out_for_next(data_out_for_next), 
		.data_in_from_next(data_in_from_next),
		.ifm_enable_write_next(ifm_enable_write_next), 
		.ifm_enable_read_next(ifm_enable_read_next), 
		.start_to_next(start_to_next)
	);
integer i,j,k;

parameter output_file = "output_file_convA2.txt";
integer output_file_id;
	initial begin
	
	output_file_id = $fopen(output_file,"w");
	
	if(!output_file_id)
	   $display("failed");
	   
		// Initialize Inputs
		clk = 0;
		reset = 1;
		riscv_data_bus = 0;
		riscv_address_bus = 0;
		data_in_from_previous = 0;
		data_in_from_next = 0;
		ifm_address_write_previous = 0;
		ifm_enable_write_previous = 0;
		start_from_previous = 0;
		end_from_next = 0;

		 
 @(negedge clk)
 reset = 0;
 

for (j=1;j<26 ; j=j+1)
begin
    for (i=2048*j; i<2048*j+1920; i=i+1)
    begin
    
    @(negedge clk)
    riscv_address_bus = i;
    riscv_data_bus =1;
    end
end

    for (k=0; k<25; k=k+1)
    begin
    @(negedge clk)
    ifm_address_write_previous = k;
    data_in_from_previous = k+1;
    ifm_enable_write_previous =1;
    end
   @(negedge clk)
   ifm_enable_write_previous = 0;
   start_from_previous = 1;
   @(negedge clk)
   start_from_previous = 0;
   
   











/*
// 1
@(negedge clk)
riscv_address_bus = 18'd2048;
riscv_data_bus = 1;

// 2
@(negedge clk)
riscv_address_bus = 18'd2049;

// 3
@(negedge clk)
riscv_address_bus = 18'd2050;

// 4
@(negedge clk)
riscv_address_bus = 18'd2051;

// 5
@(negedge clk)
riscv_address_bus = 18'd2052;
riscv_data_bus =1;

// 6
@(negedge clk)
riscv_address_bus = 18'd2053;

// memory 1
// 1
@(negedge clk)
riscv_address_bus = 18'd4096;

// 2
@(negedge clk)
riscv_address_bus = 18'd4097;
riscv_data_bus = 1;

// 4
@(negedge clk)
riscv_address_bus = 18'd4098;

// 5
@(negedge clk)
riscv_address_bus = 18'd4099;

// 6
@(negedge clk)
riscv_address_bus = 18'd4100;

// 7
@(negedge clk)
riscv_address_bus = 18'd4101;

// memory 2
// 1
@(negedge clk)
riscv_address_bus = 18'd6144;

// 2
@(negedge clk)
riscv_address_bus = 18'd6145;

// 3
@(negedge clk)
riscv_address_bus = 18'd6146;
riscv_data_bus = 1;

// 4
@(negedge clk)
riscv_address_bus = 18'd6147;

// 5
@(negedge clk)
riscv_address_bus = 18'd6148;

// 6
@(negedge clk)
riscv_address_bus = 18'd6149;

// memory 3
// 1
@(negedge clk)
riscv_address_bus = 18'd8192;

// 2
@(negedge clk)
riscv_address_bus = 18'd8193;

// 3
@(negedge clk)
riscv_address_bus = 18'd8194;

// 4
@(negedge clk)
riscv_address_bus = 18'd8195;

// 5
@(negedge clk)
riscv_address_bus = 18'd8196;
riscv_data_bus = 1;

// 6
@(negedge clk)
riscv_address_bus = 18'd8197;

// memory 4
// 1
@(negedge clk)
riscv_address_bus = 18'd10240;

// 2
@(negedge clk)
riscv_address_bus = 18'd10241;

// 3
@(negedge clk)
riscv_address_bus = 18'd10242;

// 4
@(negedge clk)
riscv_address_bus = 18'd10243;

// 5
@(negedge clk)
riscv_address_bus = 18'd10244;

// 6
@(negedge clk)
riscv_address_bus = 18'd10245;
riscv_data_bus = 1;

// memory 5
// 1
@(negedge clk)
riscv_address_bus = 18'd12288;

// 2
@(negedge clk)
riscv_address_bus = 18'd12289;

// 3
@(negedge clk)
riscv_address_bus = 18'd12290;

// 4
@(negedge clk)
riscv_address_bus = 18'd12291;

// 5
@(negedge clk)
riscv_address_bus = 18'd12292;
riscv_data_bus = 1;

// 6
@(negedge clk)
riscv_address_bus = 18'd12293;

// memory 6
// 1
@(negedge clk)
riscv_address_bus = 18'd14336;

// 2
@(negedge clk)
riscv_address_bus = 18'd14337;

// 3
@(negedge clk)
riscv_address_bus = 18'd14338;

// 4
@(negedge clk)
riscv_address_bus = 18'd14339;

// 5
@(negedge clk)
riscv_address_bus = 18'd14340;

// 6
@(negedge clk)
riscv_address_bus = 18'd14341;

// memory 7
// 1
@(negedge clk)
riscv_address_bus = 18'd16384;
riscv_data_bus = 1;

// 2
@(negedge clk)
riscv_address_bus = 18'd16385;

// 3
@(negedge clk)
riscv_address_bus = 18'd16386;

// 4
@(negedge clk)
riscv_address_bus = 18'd16387;

// 5
@(negedge clk)
riscv_address_bus = 18'd16388;

// 6
@(negedge clk)
riscv_address_bus = 18'd16389;

// memory 8
// 1
@(negedge clk)
riscv_address_bus = 18'd18432;

// 2
@(negedge clk)
riscv_address_bus = 18'd18433;

// 3
@(negedge clk)
riscv_address_bus = 18'd18434;

// 4
@(negedge clk)
riscv_address_bus = 18'd18435;

// 5
@(negedge clk)
riscv_address_bus = 18'd18436;

// 6
@(negedge clk)
riscv_address_bus = 18'd18437;

// memory 9
// 1
@(negedge clk)
riscv_address_bus = 18'd20480;

// 2
@(negedge clk)
riscv_address_bus = 18'd20481;

// 3
@(negedge clk)
riscv_address_bus = 18'd20482;

// 4
@(negedge clk)
riscv_address_bus = 18'd20483;

// 5
@(negedge clk)
riscv_address_bus = 18'd20484;

// 6
@(negedge clk)
riscv_address_bus = 18'd20485;

// memory 10
// 1
@(negedge clk)
riscv_address_bus = 18'd22528;

// 2
@(negedge clk)
riscv_address_bus = 18'd22529;

// 3
@(negedge clk)
riscv_address_bus = 18'd22530;

// 4
@(negedge clk)
riscv_address_bus = 18'd22531;

// 5
@(negedge clk)
riscv_address_bus = 18'd22532;

// 6
@(negedge clk)
riscv_address_bus = 18'd22533;

// memory 11
// 1
@(negedge clk)
riscv_address_bus = 18'd24576;

// 2
@(negedge clk)
riscv_address_bus = 18'd24577;

// 3
@(negedge clk)
riscv_address_bus = 18'd24578;

// 4
@(negedge clk)
riscv_address_bus = 18'd24579;

// 5
@(negedge clk)
riscv_address_bus = 18'd24580;

// 6
@(negedge clk)
riscv_address_bus = 18'd24581;

// memory 12
// 1
@(negedge clk)
riscv_address_bus = 18'd26624;

// 2
@(negedge clk)
riscv_address_bus = 18'd26625;

// 3
@(negedge clk)
riscv_address_bus = 18'd26626;

// 4
@(negedge clk)
riscv_address_bus = 18'd26627;

// 5
@(negedge clk)
riscv_address_bus = 18'd26628;

// 6
@(negedge clk)
riscv_address_bus = 18'd26629;

// memory 13
// 1
@(negedge clk)
riscv_address_bus = 18'd28672;

// 2
@(negedge clk)
riscv_address_bus = 18'd28673;

// 3
@(negedge clk)
riscv_address_bus = 18'd28674;

// 4
@(negedge clk)
riscv_address_bus = 18'd28675;

// 18
@(negedge clk)
riscv_address_bus = 18'd28676;

// 19
@(negedge clk)
riscv_address_bus = 18'd28677;

// memory 14
// 15
@(negedge clk)
riscv_address_bus = 18'd30720;

// 16
@(negedge clk)
riscv_address_bus = 18'd30721;

// 17
@(negedge clk)
riscv_address_bus = 18'd30722;

// 18
@(negedge clk)
riscv_address_bus = 18'd30723;

// 19
@(negedge clk)
riscv_address_bus = 18'd30724;

// 20
@(negedge clk)
riscv_address_bus = 18'd30725;

// memory 15
// 16
@(negedge clk)
riscv_address_bus = 18'd32768;

// 17
@(negedge clk)
riscv_address_bus = 18'd32769;

// 18
@(negedge clk)
riscv_address_bus = 18'd32770;

// 19
@(negedge clk)
riscv_address_bus = 18'd32771;

// 20
@(negedge clk)
riscv_address_bus = 18'd32772;

// 21
@(negedge clk)
riscv_address_bus = 18'd32773;

// memory 16
// 17
@(negedge clk)
riscv_address_bus = 18'd34816;

// 18
@(negedge clk)
riscv_address_bus = 18'd34817;

// 19
@(negedge clk)
riscv_address_bus = 18'd34818;

// 20
@(negedge clk)
riscv_address_bus = 18'd34819;

// 21
@(negedge clk)
riscv_address_bus = 18'd34820;

// 22
@(negedge clk)
riscv_address_bus = 18'd34821;

// memory 17
// 18
@(negedge clk)
riscv_address_bus = 18'd36864;

// 19
@(negedge clk)
riscv_address_bus = 18'd36865;

// 20
@(negedge clk)
riscv_address_bus = 18'd36866;

// 21
@(negedge clk)
riscv_address_bus = 18'd36867;

// 22
@(negedge clk)
riscv_address_bus = 18'd36868;

// 23
@(negedge clk)
riscv_address_bus = 18'd36869;

// memory 18
// 19
@(negedge clk)
riscv_address_bus = 18'd38912;

// 20
@(negedge clk)
riscv_address_bus = 18'd38913;

// 21
@(negedge clk)
riscv_address_bus = 18'd38914;

// 22
@(negedge clk)
riscv_address_bus = 18'd38915;

// 23
@(negedge clk)
riscv_address_bus = 18'd38916;

// 24
@(negedge clk)
riscv_address_bus = 18'd38917;

// memory 19
// 20
@(negedge clk)
riscv_address_bus = 18'd40960;

// 21
@(negedge clk)
riscv_address_bus = 18'd40961;

// 22
@(negedge clk)
riscv_address_bus = 18'd40962;

// 23
@(negedge clk)
riscv_address_bus = 18'd40963;

// 24
@(negedge clk)
riscv_address_bus = 18'd40964;

// 25
@(negedge clk)
riscv_address_bus = 18'd40965;

// memory 20
// 21
@(negedge clk)
riscv_address_bus = 18'd43008;

// 22
@(negedge clk)
riscv_address_bus = 18'd43009;

// 23
@(negedge clk)
riscv_address_bus = 18'd43010;

// 24
@(negedge clk)
riscv_address_bus = 18'd43011;

// 25
@(negedge clk)
riscv_address_bus = 18'd43012;

// 26
@(negedge clk)
riscv_address_bus = 18'd43013;

// memory 21
// 22
@(negedge clk)
riscv_address_bus = 18'd45056;

// 23
@(negedge clk)
riscv_address_bus = 18'd45057;

// 24
@(negedge clk)
riscv_address_bus = 18'd45058;

// 25
@(negedge clk)
riscv_address_bus = 18'd45059;

// 26
@(negedge clk)
riscv_address_bus = 18'd45060;

// 27
@(negedge clk)
riscv_address_bus = 18'd45061;

// memory 22
// 23
@(negedge clk)
riscv_address_bus = 18'd47104;

// 24
@(negedge clk)
riscv_address_bus = 18'd47105;

// 25
@(negedge clk)
riscv_address_bus = 18'd47106;

// 26
@(negedge clk)
riscv_address_bus = 18'd47107;

// 27
@(negedge clk)
riscv_address_bus = 18'd47108;

// 28
@(negedge clk)
riscv_address_bus = 18'd47109;

// memory 23
// 24
@(negedge clk)
riscv_address_bus = 18'd49152;

// 25
@(negedge clk)
riscv_address_bus = 18'd49153;

// 26
@(negedge clk)
riscv_address_bus = 18'd49154;

// 27
@(negedge clk)
riscv_address_bus = 18'd49155;

// 28
@(negedge clk)
riscv_address_bus = 18'd49156;

// 29
@(negedge clk)
riscv_address_bus = 18'd49157;

// memory 24
// 25
@(negedge clk)
riscv_address_bus = 18'd51200;

// 26
@(negedge clk)
riscv_address_bus = 18'd51201;

// 27
@(negedge clk)
riscv_address_bus = 18'd51202;

// 28
@(negedge clk)
riscv_address_bus = 18'd51203;

// 29
@(negedge clk)
riscv_address_bus = 18'd51204;

// 30
@(negedge clk)
riscv_address_bus = 18'd51205;

/////////////////////////////////////////
@(negedge clk)
ifm_address_write_previous = 8'd0;
ifm_enable_write_previous = 1'b1;
data_in_from_previous = 1;
@(negedge clk)
ifm_address_write_previous = 8'd1;
data_in_from_previous = 2;
@(negedge clk)
ifm_address_write_previous = 8'd2;
data_in_from_previous = 3;
@(negedge clk)
ifm_address_write_previous = 8'd3;
data_in_from_previous = 4;
@(negedge clk)
ifm_address_write_previous = 8'd4;
data_in_from_previous = 5;
@(negedge clk)
ifm_address_write_previous = 8'd5;
data_in_from_previous = 6;
@(negedge clk)
ifm_address_write_previous = 8'd6;
data_in_from_previous = 7;
@(negedge clk)
ifm_address_write_previous = 8'd7;
data_in_from_previous = 8;
@(negedge clk)
ifm_address_write_previous = 8'd8;
data_in_from_previous = 9;
@(negedge clk)
ifm_address_write_previous = 8'd9;
data_in_from_previous = 10;
@(negedge clk)
ifm_address_write_previous = 8'd10;
data_in_from_previous = 11;
@(negedge clk)
ifm_address_write_previous = 8'd11;
data_in_from_previous = 12;
@(negedge clk)
ifm_address_write_previous = 8'd12;
data_in_from_previous = 13;
@(negedge clk)
ifm_address_write_previous = 8'd13;
data_in_from_previous = 14;
@(negedge clk)
ifm_address_write_previous = 8'd14;
data_in_from_previous = 15;
@(negedge clk)
ifm_address_write_previous = 8'd15;
data_in_from_previous = 16;
@(negedge clk)
ifm_address_write_previous = 8'd16;
data_in_from_previous = 17;
@(negedge clk)
ifm_address_write_previous = 8'd17;
data_in_from_previous = 18;
@(negedge clk)
ifm_address_write_previous = 8'd18;
data_in_from_previous = 19;
@(negedge clk)
ifm_address_write_previous = 8'd19;
data_in_from_previous = 20;
@(negedge clk)
ifm_address_write_previous = 8'd20;
data_in_from_previous = 21;
@(negedge clk)
ifm_address_write_previous = 8'd21;
data_in_from_previous = 22;
@(negedge clk)
ifm_address_write_previous = 8'd22;
data_in_from_previous = 23;
@(negedge clk)
ifm_address_write_previous = 8'd23;
data_in_from_previous = 24;
@(negedge clk)
ifm_address_write_previous = 8'd24;
data_in_from_previous = 25;
@(negedge clk)
ifm_address_write_previous = 8'd25;
data_in_from_previous = 26;
@(negedge clk)
ifm_address_write_previous = 8'd26;
data_in_from_previous = 27;
@(negedge clk)
ifm_address_write_previous = 8'd27;
data_in_from_previous = 28;
@(negedge clk)
ifm_address_write_previous = 8'd28;
data_in_from_previous = 29;
@(negedge clk)
ifm_address_write_previous = 8'd29;
data_in_from_previous = 30;
@(negedge clk)
ifm_address_write_previous = 8'd30;
data_in_from_previous = 31;
@(negedge clk)
ifm_address_write_previous = 8'd31;
data_in_from_previous = 32;
@(negedge clk)
ifm_address_write_previous = 8'd32;
data_in_from_previous = 33;
@(negedge clk)
ifm_address_write_previous = 8'd33;
data_in_from_previous = 34;
@(negedge clk)
ifm_address_write_previous = 8'd34;
data_in_from_previous = 35;
@(negedge clk)
ifm_address_write_previous = 8'd35;
data_in_from_previous = 36;
@(negedge clk)
ifm_address_write_previous = 8'd36;
data_in_from_previous = 37;
@(negedge clk)
ifm_address_write_previous = 8'd37;
data_in_from_previous = 38;
@(negedge clk)
ifm_address_write_previous = 8'd38;
data_in_from_previous = 39;
@(negedge clk)
ifm_address_write_previous = 8'd39;
data_in_from_previous = 40;
@(negedge clk)
ifm_address_write_previous = 8'd40;
data_in_from_previous = 41;
@(negedge clk)
ifm_address_write_previous = 8'd41;
data_in_from_previous = 42;
@(negedge clk)
ifm_address_write_previous = 8'd42;
data_in_from_previous = 43;
@(negedge clk)
ifm_address_write_previous = 8'd43;
data_in_from_previous = 44;
@(negedge clk)
ifm_address_write_previous = 8'd44;
data_in_from_previous = 45;
@(negedge clk)
ifm_address_write_previous = 8'd45;
data_in_from_previous = 46;
@(negedge clk)
ifm_address_write_previous = 8'd46;
data_in_from_previous = 47;
@(negedge clk)
ifm_address_write_previous = 8'd47;
data_in_from_previous = 48;
@(negedge clk)
ifm_address_write_previous = 8'd48;
data_in_from_previous = 49;
@(negedge clk)
ifm_address_write_previous = 8'd49;
data_in_from_previous = 50;
@(negedge clk)
ifm_address_write_previous = 8'd50;
data_in_from_previous = 51;
@(negedge clk)
ifm_address_write_previous = 8'd51;
data_in_from_previous = 52;
@(negedge clk)
ifm_address_write_previous = 8'd52;
data_in_from_previous = 53;
@(negedge clk)
ifm_address_write_previous = 8'd53;
data_in_from_previous = 54;
@(negedge clk)
ifm_address_write_previous = 8'd54;
data_in_from_previous = 55;
@(negedge clk)
ifm_address_write_previous = 8'd55;
data_in_from_previous = 56;
@(negedge clk)
ifm_address_write_previous = 8'd56;
data_in_from_previous = 57;
@(negedge clk)
ifm_address_write_previous = 8'd57;
data_in_from_previous = 58;
@(negedge clk)
ifm_address_write_previous = 8'd58;
data_in_from_previous = 59;
@(negedge clk)
ifm_address_write_previous = 8'd59;
data_in_from_previous = 60;
@(negedge clk)
ifm_address_write_previous = 8'd60;
data_in_from_previous = 61;
@(negedge clk)
ifm_address_write_previous = 8'd61;
data_in_from_previous = 62;
@(negedge clk)
ifm_address_write_previous = 8'd62;
data_in_from_previous = 63;
@(negedge clk)
ifm_address_write_previous = 8'd63;
data_in_from_previous = 64;
@(negedge clk)
ifm_address_write_previous = 8'd64;
data_in_from_previous = 65;
@(negedge clk)
ifm_address_write_previous = 8'd65;
data_in_from_previous = 66;
@(negedge clk)
ifm_address_write_previous = 8'd66;
data_in_from_previous = 67;
@(negedge clk)
ifm_address_write_previous = 8'd67;
data_in_from_previous = 68;
@(negedge clk)
ifm_address_write_previous = 8'd68;
data_in_from_previous = 69;
@(negedge clk)
ifm_address_write_previous = 8'd69;
data_in_from_previous = 70;
@(negedge clk)
ifm_address_write_previous = 8'd70;
data_in_from_previous = 71;
@(negedge clk)
ifm_address_write_previous = 8'd71;
data_in_from_previous = 72;
@(negedge clk)
ifm_address_write_previous = 8'd72;
data_in_from_previous = 73;
@(negedge clk)
ifm_address_write_previous = 8'd73;
data_in_from_previous = 74;
@(negedge clk)
ifm_address_write_previous = 8'd74;
data_in_from_previous = 75;
@(negedge clk)
ifm_address_write_previous = 8'd75;
data_in_from_previous = 76;
@(negedge clk)
ifm_address_write_previous = 8'd76;
data_in_from_previous = 77;
@(negedge clk)
ifm_address_write_previous = 8'd77;
data_in_from_previous = 78;
@(negedge clk)
ifm_address_write_previous = 8'd78;
data_in_from_previous = 79;
@(negedge clk)
ifm_address_write_previous = 8'd79;
data_in_from_previous = 80;
@(negedge clk)
ifm_address_write_previous = 8'd80;
data_in_from_previous = 81;
@(negedge clk)
ifm_address_write_previous = 8'd81;
data_in_from_previous = 82;
@(negedge clk)
ifm_address_write_previous = 8'd82;
data_in_from_previous = 83;
@(negedge clk)
ifm_address_write_previous = 8'd83;
data_in_from_previous = 84;
@(negedge clk)
ifm_address_write_previous = 8'd84;
data_in_from_previous = 85;
@(negedge clk)
ifm_address_write_previous = 8'd85;
data_in_from_previous = 86;
@(negedge clk)
ifm_address_write_previous = 8'd86;
data_in_from_previous = 87;
@(negedge clk)
ifm_address_write_previous = 8'd87;
data_in_from_previous = 88;
@(negedge clk)
ifm_address_write_previous = 8'd88;
data_in_from_previous = 89;
@(negedge clk)
ifm_address_write_previous = 8'd89;
data_in_from_previous = 90;
@(negedge clk)
ifm_address_write_previous = 8'd90;
data_in_from_previous = 91;
@(negedge clk)
ifm_address_write_previous = 8'd91;
data_in_from_previous = 92;
@(negedge clk)
ifm_address_write_previous = 8'd92;
data_in_from_previous = 93;
@(negedge clk)
ifm_address_write_previous = 8'd93;
data_in_from_previous = 94;
@(negedge clk)
ifm_address_write_previous = 8'd94;
data_in_from_previous = 95;
@(negedge clk)
ifm_address_write_previous = 8'd95;
data_in_from_previous = 96;
@(negedge clk)
ifm_address_write_previous = 8'd96;
data_in_from_previous = 97;
@(negedge clk)
ifm_address_write_previous = 8'd97;
data_in_from_previous = 98;
@(negedge clk)
ifm_address_write_previous = 8'd98;
data_in_from_previous = 99;
@(negedge clk)
ifm_address_write_previous = 8'd99;
data_in_from_previous = 100;
@(negedge clk)
ifm_address_write_previous = 8'd100;
data_in_from_previous = 101;
@(negedge clk)
ifm_address_write_previous = 8'd101;
data_in_from_previous = 102;
@(negedge clk)
ifm_address_write_previous = 8'd102;
data_in_from_previous = 103;
@(negedge clk)
ifm_address_write_previous = 8'd103;
data_in_from_previous = 104;
@(negedge clk)
ifm_address_write_previous = 8'd104;
data_in_from_previous = 105;
@(negedge clk)
ifm_address_write_previous = 8'd105;
data_in_from_previous = 106;
@(negedge clk)
ifm_address_write_previous = 8'd106;
data_in_from_previous = 107;
@(negedge clk)
ifm_address_write_previous = 8'd107;
data_in_from_previous = 108;
@(negedge clk)
ifm_address_write_previous = 8'd108;
data_in_from_previous = 109;
@(negedge clk)
ifm_address_write_previous = 8'd109;
data_in_from_previous = 110;
@(negedge clk)
ifm_address_write_previous = 8'd110;
data_in_from_previous = 111;
@(negedge clk)
ifm_address_write_previous = 8'd111;
data_in_from_previous = 112;
@(negedge clk)
ifm_address_write_previous = 8'd112;
data_in_from_previous = 113;
@(negedge clk)
ifm_address_write_previous = 8'd113;
data_in_from_previous = 114;
@(negedge clk)
ifm_address_write_previous = 8'd114;
data_in_from_previous = 115;
@(negedge clk)
ifm_address_write_previous = 8'd115;
data_in_from_previous = 116;
@(negedge clk)
ifm_address_write_previous = 8'd116;
data_in_from_previous = 117;
@(negedge clk)
ifm_address_write_previous = 8'd117;
data_in_from_previous = 118;
@(negedge clk)
ifm_address_write_previous = 8'd118;
data_in_from_previous = 119;
@(negedge clk)
ifm_address_write_previous = 8'd119;
data_in_from_previous = 120;
@(negedge clk)
ifm_address_write_previous = 8'd120;
data_in_from_previous = 121;
@(negedge clk)
ifm_address_write_previous = 8'd121;
data_in_from_previous = 122;
@(negedge clk)
ifm_address_write_previous = 8'd122;
data_in_from_previous = 123;
@(negedge clk)
ifm_address_write_previous = 8'd123;
data_in_from_previous = 124;
@(negedge clk)
ifm_address_write_previous = 8'd124;
data_in_from_previous = 125;
@(negedge clk)
ifm_address_write_previous = 8'd125;
data_in_from_previous = 126;
@(negedge clk)
ifm_address_write_previous = 8'd126;
data_in_from_previous = 127;
@(negedge clk)
ifm_address_write_previous = 8'd127;
data_in_from_previous = 128;
@(negedge clk)
ifm_address_write_previous = 8'd128;
data_in_from_previous = 129;
@(negedge clk)
ifm_address_write_previous = 8'd129;
data_in_from_previous = 130;
@(negedge clk)
ifm_address_write_previous = 8'd130;
data_in_from_previous = 131;
@(negedge clk)
ifm_address_write_previous = 8'd131;
data_in_from_previous = 132;
@(negedge clk)
ifm_address_write_previous = 8'd132;
data_in_from_previous = 133;
@(negedge clk)
ifm_address_write_previous = 8'd133;
data_in_from_previous = 134;
@(negedge clk)
ifm_address_write_previous = 8'd134;
data_in_from_previous = 135;
@(negedge clk)
ifm_address_write_previous = 8'd135;
data_in_from_previous = 136;
@(negedge clk)
ifm_address_write_previous = 8'd136;
data_in_from_previous = 137;
@(negedge clk)
ifm_address_write_previous = 8'd137;
data_in_from_previous = 138;
@(negedge clk)
ifm_address_write_previous = 8'd138;
data_in_from_previous = 139;
@(negedge clk)
ifm_address_write_previous = 8'd139;
data_in_from_previous = 140;
@(negedge clk)
ifm_address_write_previous = 8'd140;
data_in_from_previous = 141;
@(negedge clk)
ifm_address_write_previous = 8'd141;
data_in_from_previous = 142;
@(negedge clk)
ifm_address_write_previous = 8'd142;
data_in_from_previous = 143;
@(negedge clk)
ifm_address_write_previous = 8'd143;
data_in_from_previous = 144;
@(negedge clk)
ifm_address_write_previous = 8'd144;
data_in_from_previous = 145;
@(negedge clk)
ifm_address_write_previous = 8'd145;
data_in_from_previous = 146;
@(negedge clk)
ifm_address_write_previous = 8'd146;
data_in_from_previous = 147;
@(negedge clk)
ifm_address_write_previous = 8'd147;
data_in_from_previous = 148;
@(negedge clk)
ifm_address_write_previous = 8'd148;
data_in_from_previous = 149;
@(negedge clk)
ifm_address_write_previous = 8'd149;
data_in_from_previous = 150;
@(negedge clk)
ifm_address_write_previous = 8'd150;
data_in_from_previous = 151;
@(negedge clk)
ifm_address_write_previous = 8'd151;
data_in_from_previous = 152;
@(negedge clk)
ifm_address_write_previous = 8'd152;
data_in_from_previous = 153;
@(negedge clk)
ifm_address_write_previous = 8'd153;
data_in_from_previous = 154;
@(negedge clk)
ifm_address_write_previous = 8'd154;
data_in_from_previous = 155;
@(negedge clk)
ifm_address_write_previous = 8'd155;
data_in_from_previous = 156;
@(negedge clk)
ifm_address_write_previous = 8'd156;
data_in_from_previous = 157;
@(negedge clk)
ifm_address_write_previous = 8'd157;
data_in_from_previous = 158;
@(negedge clk)
ifm_address_write_previous = 8'd158;
data_in_from_previous = 159;
@(negedge clk)
ifm_address_write_previous = 8'd159;
data_in_from_previous = 160;
@(negedge clk)
ifm_address_write_previous = 8'd160;
data_in_from_previous = 161;
@(negedge clk)
ifm_address_write_previous = 8'd161;
data_in_from_previous = 162;
@(negedge clk)
ifm_address_write_previous = 8'd162;
data_in_from_previous = 163;
@(negedge clk)
ifm_address_write_previous = 8'd163;
data_in_from_previous = 164;
@(negedge clk)
ifm_address_write_previous = 8'd164;
data_in_from_previous = 165;
@(negedge clk)
ifm_address_write_previous = 8'd165;
data_in_from_previous = 166;
@(negedge clk)
ifm_address_write_previous = 8'd166;
data_in_from_previous = 167;
@(negedge clk)
ifm_address_write_previous = 8'd167;
data_in_from_previous = 168;
@(negedge clk)
ifm_address_write_previous = 8'd168;
data_in_from_previous = 169;
@(negedge clk)
ifm_address_write_previous = 8'd169;
data_in_from_previous = 170;
@(negedge clk)
ifm_address_write_previous = 8'd170;
data_in_from_previous = 171;
@(negedge clk)
ifm_address_write_previous = 8'd171;
data_in_from_previous = 172;
@(negedge clk)
ifm_address_write_previous = 8'd172;
data_in_from_previous = 173;
@(negedge clk)
ifm_address_write_previous = 8'd173;
data_in_from_previous = 174;
@(negedge clk)
ifm_address_write_previous = 8'd174;
data_in_from_previous = 175;
@(negedge clk)
ifm_address_write_previous = 8'd175;
data_in_from_previous = 176;
@(negedge clk)
ifm_address_write_previous = 8'd176;
data_in_from_previous = 177;
@(negedge clk)
ifm_address_write_previous = 8'd177;
data_in_from_previous = 178;
@(negedge clk)
ifm_address_write_previous = 8'd178;
data_in_from_previous = 179;
@(negedge clk)
ifm_address_write_previous = 8'd179;
data_in_from_previous = 180;
@(negedge clk)
ifm_address_write_previous = 8'd180;
data_in_from_previous = 181;
@(negedge clk)
ifm_address_write_previous = 8'd181;
data_in_from_previous = 182;
@(negedge clk)
ifm_address_write_previous = 8'd182;
data_in_from_previous = 183;
@(negedge clk)
ifm_address_write_previous = 8'd183;
data_in_from_previous = 184;
@(negedge clk)
ifm_address_write_previous = 8'd184;
data_in_from_previous = 185;
@(negedge clk)
ifm_address_write_previous = 8'd185;
data_in_from_previous = 186;
@(negedge clk)
ifm_address_write_previous = 8'd186;
data_in_from_previous = 187;
@(negedge clk)
ifm_address_write_previous = 8'd187;
data_in_from_previous = 188;
@(negedge clk)
ifm_address_write_previous = 8'd188;
data_in_from_previous = 189;
@(negedge clk)
ifm_address_write_previous = 8'd189;
data_in_from_previous = 190;
@(negedge clk)
ifm_address_write_previous = 8'd190;
data_in_from_previous = 191;
@(negedge clk)
ifm_address_write_previous = 8'd191;
data_in_from_previous = 192;
@(negedge clk)
ifm_address_write_previous = 8'd192;
data_in_from_previous = 193;
@(negedge clk)
ifm_address_write_previous = 8'd193;
data_in_from_previous = 194;
@(negedge clk)
ifm_address_write_previous = 8'd194;
data_in_from_previous = 195;
@(negedge clk)
ifm_address_write_previous = 8'd195;
data_in_from_previous = 196;
@(negedge clk)
start_from_previous = 1'b1;
ifm_enable_write_previous = 1'b0;
@(negedge clk)
start_from_previous = 1'b0;
@(negedge clk)
ifm_address_write_previous = 8'd0;
ifm_enable_write_previous = 1'b1;
data_in_from_previous = 1;
@(negedge clk)
ifm_address_write_previous = 8'd1;
data_in_from_previous = 2;
@(negedge clk)
ifm_address_write_previous = 8'd2;
data_in_from_previous = 3;
@(negedge clk)
ifm_address_write_previous = 8'd3;
data_in_from_previous = 4;
@(negedge clk)
ifm_address_write_previous = 8'd4;
data_in_from_previous = 5;
@(negedge clk)
ifm_address_write_previous = 8'd5;
data_in_from_previous = 6;
@(negedge clk)
ifm_address_write_previous = 8'd6;
data_in_from_previous = 7;
@(negedge clk)
ifm_address_write_previous = 8'd7;
data_in_from_previous = 8;
@(negedge clk)
ifm_address_write_previous = 8'd8;
data_in_from_previous = 9;
@(negedge clk)
ifm_address_write_previous = 8'd9;
data_in_from_previous = 10;
@(negedge clk)
ifm_address_write_previous = 8'd10;
data_in_from_previous = 11;
@(negedge clk)
ifm_address_write_previous = 8'd11;
data_in_from_previous = 12;
@(negedge clk)
ifm_address_write_previous = 8'd12;
data_in_from_previous = 13;
@(negedge clk)
ifm_address_write_previous = 8'd13;
data_in_from_previous = 14;
@(negedge clk)
ifm_address_write_previous = 8'd14;
data_in_from_previous = 15;
@(negedge clk)
ifm_address_write_previous = 8'd15;
data_in_from_previous = 16;
@(negedge clk)
ifm_address_write_previous = 8'd16;
data_in_from_previous = 17;
@(negedge clk)
ifm_address_write_previous = 8'd17;
data_in_from_previous = 18;
@(negedge clk)
ifm_address_write_previous = 8'd18;
data_in_from_previous = 19;
@(negedge clk)
ifm_address_write_previous = 8'd19;
data_in_from_previous = 20;
@(negedge clk)
ifm_address_write_previous = 8'd20;
data_in_from_previous = 21;
@(negedge clk)
ifm_address_write_previous = 8'd21;
data_in_from_previous = 22;
@(negedge clk)
ifm_address_write_previous = 8'd22;
data_in_from_previous = 23;
@(negedge clk)
ifm_address_write_previous = 8'd23;
data_in_from_previous = 24;
@(negedge clk)
ifm_address_write_previous = 8'd24;
data_in_from_previous = 25;
@(negedge clk)
ifm_address_write_previous = 8'd25;
data_in_from_previous = 26;
@(negedge clk)
ifm_address_write_previous = 8'd26;
data_in_from_previous = 27;
@(negedge clk)
ifm_address_write_previous = 8'd27;
data_in_from_previous = 28;
@(negedge clk)
ifm_address_write_previous = 8'd28;
data_in_from_previous = 29;
@(negedge clk)
ifm_address_write_previous = 8'd29;
data_in_from_previous = 30;
@(negedge clk)
ifm_address_write_previous = 8'd30;
data_in_from_previous = 31;
@(negedge clk)
ifm_address_write_previous = 8'd31;
data_in_from_previous = 32;
@(negedge clk)
ifm_address_write_previous = 8'd32;
data_in_from_previous = 33;
@(negedge clk)
ifm_address_write_previous = 8'd33;
data_in_from_previous = 34;
@(negedge clk)
ifm_address_write_previous = 8'd34;
data_in_from_previous = 35;
@(negedge clk)
ifm_address_write_previous = 8'd35;
data_in_from_previous = 36;
@(negedge clk)
ifm_address_write_previous = 8'd36;
data_in_from_previous = 37;
@(negedge clk)
ifm_address_write_previous = 8'd37;
data_in_from_previous = 38;
@(negedge clk)
ifm_address_write_previous = 8'd38;
data_in_from_previous = 39;
@(negedge clk)
ifm_address_write_previous = 8'd39;
data_in_from_previous = 40;
@(negedge clk)
ifm_address_write_previous = 8'd40;
data_in_from_previous = 41;
@(negedge clk)
ifm_address_write_previous = 8'd41;
data_in_from_previous = 42;
@(negedge clk)
ifm_address_write_previous = 8'd42;
data_in_from_previous = 43;
@(negedge clk)
ifm_address_write_previous = 8'd43;
data_in_from_previous = 44;
@(negedge clk)
ifm_address_write_previous = 8'd44;
data_in_from_previous = 45;
@(negedge clk)
ifm_address_write_previous = 8'd45;
data_in_from_previous = 46;
@(negedge clk)
ifm_address_write_previous = 8'd46;
data_in_from_previous = 47;
@(negedge clk)
ifm_address_write_previous = 8'd47;
data_in_from_previous = 48;
@(negedge clk)
ifm_address_write_previous = 8'd48;
data_in_from_previous = 49;
@(negedge clk)
ifm_address_write_previous = 8'd49;
data_in_from_previous = 50;
@(negedge clk)
ifm_address_write_previous = 8'd50;
data_in_from_previous = 51;
@(negedge clk)
ifm_address_write_previous = 8'd51;
data_in_from_previous = 52;
@(negedge clk)
ifm_address_write_previous = 8'd52;
data_in_from_previous = 53;
@(negedge clk)
ifm_address_write_previous = 8'd53;
data_in_from_previous = 54;
@(negedge clk)
ifm_address_write_previous = 8'd54;
data_in_from_previous = 55;
@(negedge clk)
ifm_address_write_previous = 8'd55;
data_in_from_previous = 56;
@(negedge clk)
ifm_address_write_previous = 8'd56;
data_in_from_previous = 57;
@(negedge clk)
ifm_address_write_previous = 8'd57;
data_in_from_previous = 58;
@(negedge clk)
ifm_address_write_previous = 8'd58;
data_in_from_previous = 59;
@(negedge clk)
ifm_address_write_previous = 8'd59;
data_in_from_previous = 60;
@(negedge clk)
ifm_address_write_previous = 8'd60;
data_in_from_previous = 61;
@(negedge clk)
ifm_address_write_previous = 8'd61;
data_in_from_previous = 62;
@(negedge clk)
ifm_address_write_previous = 8'd62;
data_in_from_previous = 63;
@(negedge clk)
ifm_address_write_previous = 8'd63;
data_in_from_previous = 64;
@(negedge clk)
ifm_address_write_previous = 8'd64;
data_in_from_previous = 65;
@(negedge clk)
ifm_address_write_previous = 8'd65;
data_in_from_previous = 66;
@(negedge clk)
ifm_address_write_previous = 8'd66;
data_in_from_previous = 67;
@(negedge clk)
ifm_address_write_previous = 8'd67;
data_in_from_previous = 68;
@(negedge clk)
ifm_address_write_previous = 8'd68;
data_in_from_previous = 69;
@(negedge clk)
ifm_address_write_previous = 8'd69;
data_in_from_previous = 70;
@(negedge clk)
ifm_address_write_previous = 8'd70;
data_in_from_previous = 71;
@(negedge clk)
ifm_address_write_previous = 8'd71;
data_in_from_previous = 72;
@(negedge clk)
ifm_address_write_previous = 8'd72;
data_in_from_previous = 73;
@(negedge clk)
ifm_address_write_previous = 8'd73;
data_in_from_previous = 74;
@(negedge clk)
ifm_address_write_previous = 8'd74;
data_in_from_previous = 75;
@(negedge clk)
ifm_address_write_previous = 8'd75;
data_in_from_previous = 76;
@(negedge clk)
ifm_address_write_previous = 8'd76;
data_in_from_previous = 77;
@(negedge clk)
ifm_address_write_previous = 8'd77;
data_in_from_previous = 78;
@(negedge clk)
ifm_address_write_previous = 8'd78;
data_in_from_previous = 79;
@(negedge clk)
ifm_address_write_previous = 8'd79;
data_in_from_previous = 80;
@(negedge clk)
ifm_address_write_previous = 8'd80;
data_in_from_previous = 81;
@(negedge clk)
ifm_address_write_previous = 8'd81;
data_in_from_previous = 82;
@(negedge clk)
ifm_address_write_previous = 8'd82;
data_in_from_previous = 83;
@(negedge clk)
ifm_address_write_previous = 8'd83;
data_in_from_previous = 84;
@(negedge clk)
ifm_address_write_previous = 8'd84;
data_in_from_previous = 85;
@(negedge clk)
ifm_address_write_previous = 8'd85;
data_in_from_previous = 86;
@(negedge clk)
ifm_address_write_previous = 8'd86;
data_in_from_previous = 87;
@(negedge clk)
ifm_address_write_previous = 8'd87;
data_in_from_previous = 88;
@(negedge clk)
ifm_address_write_previous = 8'd88;
data_in_from_previous = 89;
@(negedge clk)
ifm_address_write_previous = 8'd89;
data_in_from_previous = 90;
@(negedge clk)
ifm_address_write_previous = 8'd90;
data_in_from_previous = 91;
@(negedge clk)
ifm_address_write_previous = 8'd91;
data_in_from_previous = 92;
@(negedge clk)
ifm_address_write_previous = 8'd92;
data_in_from_previous = 93;
@(negedge clk)
ifm_address_write_previous = 8'd93;
data_in_from_previous = 94;
@(negedge clk)
ifm_address_write_previous = 8'd94;
data_in_from_previous = 95;
@(negedge clk)
ifm_address_write_previous = 8'd95;
data_in_from_previous = 96;
@(negedge clk)
ifm_address_write_previous = 8'd96;
data_in_from_previous = 97;
@(negedge clk)
ifm_address_write_previous = 8'd97;
data_in_from_previous = 98;
@(negedge clk)
ifm_address_write_previous = 8'd98;
data_in_from_previous = 99;
@(negedge clk)
ifm_address_write_previous = 8'd99;
data_in_from_previous = 100;
@(negedge clk)
ifm_address_write_previous = 8'd100;
data_in_from_previous = 101;
@(negedge clk)
ifm_address_write_previous = 8'd101;
data_in_from_previous = 102;
@(negedge clk)
ifm_address_write_previous = 8'd102;
data_in_from_previous = 103;
@(negedge clk)
ifm_address_write_previous = 8'd103;
data_in_from_previous = 104;
@(negedge clk)
ifm_address_write_previous = 8'd104;
data_in_from_previous = 105;
@(negedge clk)
ifm_address_write_previous = 8'd105;
data_in_from_previous = 106;
@(negedge clk)
ifm_address_write_previous = 8'd106;
data_in_from_previous = 107;
@(negedge clk)
ifm_address_write_previous = 8'd107;
data_in_from_previous = 108;
@(negedge clk)
ifm_address_write_previous = 8'd108;
data_in_from_previous = 109;
@(negedge clk)
ifm_address_write_previous = 8'd109;
data_in_from_previous = 110;
@(negedge clk)
ifm_address_write_previous = 8'd110;
data_in_from_previous = 111;
@(negedge clk)
ifm_address_write_previous = 8'd111;
data_in_from_previous = 112;
@(negedge clk)
ifm_address_write_previous = 8'd112;
data_in_from_previous = 113;
@(negedge clk)
ifm_address_write_previous = 8'd113;
data_in_from_previous = 114;
@(negedge clk)
ifm_address_write_previous = 8'd114;
data_in_from_previous = 115;
@(negedge clk)
ifm_address_write_previous = 8'd115;
data_in_from_previous = 116;
@(negedge clk)
ifm_address_write_previous = 8'd116;
data_in_from_previous = 117;
@(negedge clk)
ifm_address_write_previous = 8'd117;
data_in_from_previous = 118;
@(negedge clk)
ifm_address_write_previous = 8'd118;
data_in_from_previous = 119;
@(negedge clk)
ifm_address_write_previous = 8'd119;
data_in_from_previous = 120;
@(negedge clk)
ifm_address_write_previous = 8'd120;
data_in_from_previous = 121;
@(negedge clk)
ifm_address_write_previous = 8'd121;
data_in_from_previous = 122;
@(negedge clk)
ifm_address_write_previous = 8'd122;
data_in_from_previous = 123;
@(negedge clk)
ifm_address_write_previous = 8'd123;
data_in_from_previous = 124;
@(negedge clk)
ifm_address_write_previous = 8'd124;
data_in_from_previous = 125;
@(negedge clk)
ifm_address_write_previous = 8'd125;
data_in_from_previous = 126;
@(negedge clk)
ifm_address_write_previous = 8'd126;
data_in_from_previous = 127;
@(negedge clk)
ifm_address_write_previous = 8'd127;
data_in_from_previous = 128;
@(negedge clk)
ifm_address_write_previous = 8'd128;
data_in_from_previous = 129;
@(negedge clk)
ifm_address_write_previous = 8'd129;
data_in_from_previous = 130;
@(negedge clk)
ifm_address_write_previous = 8'd130;
data_in_from_previous = 131;
@(negedge clk)
ifm_address_write_previous = 8'd131;
data_in_from_previous = 132;
@(negedge clk)
ifm_address_write_previous = 8'd132;
data_in_from_previous = 133;
@(negedge clk)
ifm_address_write_previous = 8'd133;
data_in_from_previous = 134;
@(negedge clk)
ifm_address_write_previous = 8'd134;
data_in_from_previous = 135;
@(negedge clk)
ifm_address_write_previous = 8'd135;
data_in_from_previous = 136;
@(negedge clk)
ifm_address_write_previous = 8'd136;
data_in_from_previous = 137;
@(negedge clk)
ifm_address_write_previous = 8'd137;
data_in_from_previous = 138;
@(negedge clk)
ifm_address_write_previous = 8'd138;
data_in_from_previous = 139;
@(negedge clk)
ifm_address_write_previous = 8'd139;
data_in_from_previous = 140;
@(negedge clk)
ifm_address_write_previous = 8'd140;
data_in_from_previous = 141;
@(negedge clk)
ifm_address_write_previous = 8'd141;
data_in_from_previous = 142;
@(negedge clk)
ifm_address_write_previous = 8'd142;
data_in_from_previous = 143;
@(negedge clk)
ifm_address_write_previous = 8'd143;
data_in_from_previous = 144;
@(negedge clk)
ifm_address_write_previous = 8'd144;
data_in_from_previous = 145;
@(negedge clk)
ifm_address_write_previous = 8'd145;
data_in_from_previous = 146;
@(negedge clk)
ifm_address_write_previous = 8'd146;
data_in_from_previous = 147;
@(negedge clk)
ifm_address_write_previous = 8'd147;
data_in_from_previous = 148;
@(negedge clk)
ifm_address_write_previous = 8'd148;
data_in_from_previous = 149;
@(negedge clk)
ifm_address_write_previous = 8'd149;
data_in_from_previous = 150;
@(negedge clk)
ifm_address_write_previous = 8'd150;
data_in_from_previous = 151;
@(negedge clk)
ifm_address_write_previous = 8'd151;
data_in_from_previous = 152;
@(negedge clk)
ifm_address_write_previous = 8'd152;
data_in_from_previous = 153;
@(negedge clk)
ifm_address_write_previous = 8'd153;
data_in_from_previous = 154;
@(negedge clk)
ifm_address_write_previous = 8'd154;
data_in_from_previous = 155;
@(negedge clk)
ifm_address_write_previous = 8'd155;
data_in_from_previous = 156;
@(negedge clk)
ifm_address_write_previous = 8'd156;
data_in_from_previous = 157;
@(negedge clk)
ifm_address_write_previous = 8'd157;
data_in_from_previous = 158;
@(negedge clk)
ifm_address_write_previous = 8'd158;
data_in_from_previous = 159;
@(negedge clk)
ifm_address_write_previous = 8'd159;
data_in_from_previous = 160;
@(negedge clk)
ifm_address_write_previous = 8'd160;
data_in_from_previous = 161;
@(negedge clk)
ifm_address_write_previous = 8'd161;
data_in_from_previous = 162;
@(negedge clk)
ifm_address_write_previous = 8'd162;
data_in_from_previous = 163;
@(negedge clk)
ifm_address_write_previous = 8'd163;
data_in_from_previous = 164;
@(negedge clk)
ifm_address_write_previous = 8'd164;
data_in_from_previous = 165;
@(negedge clk)
ifm_address_write_previous = 8'd165;
data_in_from_previous = 166;
@(negedge clk)
ifm_address_write_previous = 8'd166;
data_in_from_previous = 167;
@(negedge clk)
ifm_address_write_previous = 8'd167;
data_in_from_previous = 168;
@(negedge clk)
ifm_address_write_previous = 8'd168;
data_in_from_previous = 169;
@(negedge clk)
ifm_address_write_previous = 8'd169;
data_in_from_previous = 170;
@(negedge clk)
ifm_address_write_previous = 8'd170;
data_in_from_previous = 171;
@(negedge clk)
ifm_address_write_previous = 8'd171;
data_in_from_previous = 172;
@(negedge clk)
ifm_address_write_previous = 8'd172;
data_in_from_previous = 173;
@(negedge clk)
ifm_address_write_previous = 8'd173;
data_in_from_previous = 174;
@(negedge clk)
ifm_address_write_previous = 8'd174;
data_in_from_previous = 175;
@(negedge clk)
ifm_address_write_previous = 8'd175;
data_in_from_previous = 176;
@(negedge clk)
ifm_address_write_previous = 8'd176;
data_in_from_previous = 177;
@(negedge clk)
ifm_address_write_previous = 8'd177;
data_in_from_previous = 178;
@(negedge clk)
ifm_address_write_previous = 8'd178;
data_in_from_previous = 179;
@(negedge clk)
ifm_address_write_previous = 8'd179;
data_in_from_previous = 180;
@(negedge clk)
ifm_address_write_previous = 8'd180;
data_in_from_previous = 181;
@(negedge clk)
ifm_address_write_previous = 8'd181;
data_in_from_previous = 182;
@(negedge clk)
ifm_address_write_previous = 8'd182;
data_in_from_previous = 183;
@(negedge clk)
ifm_address_write_previous = 8'd183;
data_in_from_previous = 184;
@(negedge clk)
ifm_address_write_previous = 8'd184;
data_in_from_previous = 185;
@(negedge clk)
ifm_address_write_previous = 8'd185;
data_in_from_previous = 186;
@(negedge clk)
ifm_address_write_previous = 8'd186;
data_in_from_previous = 187;
@(negedge clk)
ifm_address_write_previous = 8'd187;
data_in_from_previous = 188;
@(negedge clk)
ifm_address_write_previous = 8'd188;
data_in_from_previous = 189;
@(negedge clk)
ifm_address_write_previous = 8'd189;
data_in_from_previous = 190;
@(negedge clk)
ifm_address_write_previous = 8'd190;
data_in_from_previous = 191;
@(negedge clk)
ifm_address_write_previous = 8'd191;
data_in_from_previous = 192;
@(negedge clk)
ifm_address_write_previous = 8'd192;
data_in_from_previous = 193;
@(negedge clk)
ifm_address_write_previous = 8'd193;
data_in_from_previous = 194;
@(negedge clk)
ifm_address_write_previous = 8'd194;
data_in_from_previous = 195;
@(negedge clk)
ifm_address_write_previous = 8'd195;
data_in_from_previous = 196;
@(negedge clk)
ifm_enable_write_previous = 1'b0;
#13900
@(negedge clk)
start_from_previous = 1'b1;
ifm_enable_write_previous = 1'b0;
@(negedge clk)
start_from_previous = 1'b0;
@(negedge clk)
ifm_address_write_previous = 8'd0;
ifm_enable_write_previous = 1'b1;
data_in_from_previous = 1;
@(negedge clk)
ifm_address_write_previous = 8'd1;
data_in_from_previous = 2;
@(negedge clk)
ifm_address_write_previous = 8'd2;
data_in_from_previous = 3;
@(negedge clk)
ifm_address_write_previous = 8'd3;
data_in_from_previous = 4;
@(negedge clk)
ifm_address_write_previous = 8'd4;
data_in_from_previous = 5;
@(negedge clk)
ifm_address_write_previous = 8'd5;
data_in_from_previous = 6;
@(negedge clk)
ifm_address_write_previous = 8'd6;
data_in_from_previous = 7;
@(negedge clk)
ifm_address_write_previous = 8'd7;
data_in_from_previous = 8;
@(negedge clk)
ifm_address_write_previous = 8'd8;
data_in_from_previous = 9;
@(negedge clk)
ifm_address_write_previous = 8'd9;
data_in_from_previous = 10;
@(negedge clk)
ifm_address_write_previous = 8'd10;
data_in_from_previous = 11;
@(negedge clk)
ifm_address_write_previous = 8'd11;
data_in_from_previous = 12;
@(negedge clk)
ifm_address_write_previous = 8'd12;
data_in_from_previous = 13;
@(negedge clk)
ifm_address_write_previous = 8'd13;
data_in_from_previous = 14;
@(negedge clk)
ifm_address_write_previous = 8'd14;
data_in_from_previous = 15;
@(negedge clk)
ifm_address_write_previous = 8'd15;
data_in_from_previous = 16;
@(negedge clk)
ifm_address_write_previous = 8'd16;
data_in_from_previous = 17;
@(negedge clk)
ifm_address_write_previous = 8'd17;
data_in_from_previous = 18;
@(negedge clk)
ifm_address_write_previous = 8'd18;
data_in_from_previous = 19;
@(negedge clk)
ifm_address_write_previous = 8'd19;
data_in_from_previous = 20;
@(negedge clk)
ifm_address_write_previous = 8'd20;
data_in_from_previous = 21;
@(negedge clk)
ifm_address_write_previous = 8'd21;
data_in_from_previous = 22;
@(negedge clk)
ifm_address_write_previous = 8'd22;
data_in_from_previous = 23;
@(negedge clk)
ifm_address_write_previous = 8'd23;
data_in_from_previous = 24;
@(negedge clk)
ifm_address_write_previous = 8'd24;
data_in_from_previous = 25;
@(negedge clk)
ifm_address_write_previous = 8'd25;
data_in_from_previous = 26;
@(negedge clk)
ifm_address_write_previous = 8'd26;
data_in_from_previous = 27;
@(negedge clk)
ifm_address_write_previous = 8'd27;
data_in_from_previous = 28;
@(negedge clk)
ifm_address_write_previous = 8'd28;
data_in_from_previous = 29;
@(negedge clk)
ifm_address_write_previous = 8'd29;
data_in_from_previous = 30;
@(negedge clk)
ifm_address_write_previous = 8'd30;
data_in_from_previous = 31;
@(negedge clk)
ifm_address_write_previous = 8'd31;
data_in_from_previous = 32;
@(negedge clk)
ifm_address_write_previous = 8'd32;
data_in_from_previous = 33;
@(negedge clk)
ifm_address_write_previous = 8'd33;
data_in_from_previous = 34;
@(negedge clk)
ifm_address_write_previous = 8'd34;
data_in_from_previous = 35;
@(negedge clk)
ifm_address_write_previous = 8'd35;
data_in_from_previous = 36;
@(negedge clk)
ifm_address_write_previous = 8'd36;
data_in_from_previous = 37;
@(negedge clk)
ifm_address_write_previous = 8'd37;
data_in_from_previous = 38;
@(negedge clk)
ifm_address_write_previous = 8'd38;
data_in_from_previous = 39;
@(negedge clk)
ifm_address_write_previous = 8'd39;
data_in_from_previous = 40;
@(negedge clk)
ifm_address_write_previous = 8'd40;
data_in_from_previous = 41;
@(negedge clk)
ifm_address_write_previous = 8'd41;
data_in_from_previous = 42;
@(negedge clk)
ifm_address_write_previous = 8'd42;
data_in_from_previous = 43;
@(negedge clk)
ifm_address_write_previous = 8'd43;
data_in_from_previous = 44;
@(negedge clk)
ifm_address_write_previous = 8'd44;
data_in_from_previous = 45;
@(negedge clk)
ifm_address_write_previous = 8'd45;
data_in_from_previous = 46;
@(negedge clk)
ifm_address_write_previous = 8'd46;
data_in_from_previous = 47;
@(negedge clk)
ifm_address_write_previous = 8'd47;
data_in_from_previous = 48;
@(negedge clk)
ifm_address_write_previous = 8'd48;
data_in_from_previous = 49;
@(negedge clk)
ifm_address_write_previous = 8'd49;
data_in_from_previous = 50;
@(negedge clk)
ifm_address_write_previous = 8'd50;
data_in_from_previous = 51;
@(negedge clk)
ifm_address_write_previous = 8'd51;
data_in_from_previous = 52;
@(negedge clk)
ifm_address_write_previous = 8'd52;
data_in_from_previous = 53;
@(negedge clk)
ifm_address_write_previous = 8'd53;
data_in_from_previous = 54;
@(negedge clk)
ifm_address_write_previous = 8'd54;
data_in_from_previous = 55;
@(negedge clk)
ifm_address_write_previous = 8'd55;
data_in_from_previous = 56;
@(negedge clk)
ifm_address_write_previous = 8'd56;
data_in_from_previous = 57;
@(negedge clk)
ifm_address_write_previous = 8'd57;
data_in_from_previous = 58;
@(negedge clk)
ifm_address_write_previous = 8'd58;
data_in_from_previous = 59;
@(negedge clk)
ifm_address_write_previous = 8'd59;
data_in_from_previous = 60;
@(negedge clk)
ifm_address_write_previous = 8'd60;
data_in_from_previous = 61;
@(negedge clk)
ifm_address_write_previous = 8'd61;
data_in_from_previous = 62;
@(negedge clk)
ifm_address_write_previous = 8'd62;
data_in_from_previous = 63;
@(negedge clk)
ifm_address_write_previous = 8'd63;
data_in_from_previous = 64;
@(negedge clk)
ifm_address_write_previous = 8'd64;
data_in_from_previous = 65;
@(negedge clk)
ifm_address_write_previous = 8'd65;
data_in_from_previous = 66;
@(negedge clk)
ifm_address_write_previous = 8'd66;
data_in_from_previous = 67;
@(negedge clk)
ifm_address_write_previous = 8'd67;
data_in_from_previous = 68;
@(negedge clk)
ifm_address_write_previous = 8'd68;
data_in_from_previous = 69;
@(negedge clk)
ifm_address_write_previous = 8'd69;
data_in_from_previous = 70;
@(negedge clk)
ifm_address_write_previous = 8'd70;
data_in_from_previous = 71;
@(negedge clk)
ifm_address_write_previous = 8'd71;
data_in_from_previous = 72;
@(negedge clk)
ifm_address_write_previous = 8'd72;
data_in_from_previous = 73;
@(negedge clk)
ifm_address_write_previous = 8'd73;
data_in_from_previous = 74;
@(negedge clk)
ifm_address_write_previous = 8'd74;
data_in_from_previous = 75;
@(negedge clk)
ifm_address_write_previous = 8'd75;
data_in_from_previous = 76;
@(negedge clk)
ifm_address_write_previous = 8'd76;
data_in_from_previous = 77;
@(negedge clk)
ifm_address_write_previous = 8'd77;
data_in_from_previous = 78;
@(negedge clk)
ifm_address_write_previous = 8'd78;
data_in_from_previous = 79;
@(negedge clk)
ifm_address_write_previous = 8'd79;
data_in_from_previous = 80;
@(negedge clk)
ifm_address_write_previous = 8'd80;
data_in_from_previous = 81;
@(negedge clk)
ifm_address_write_previous = 8'd81;
data_in_from_previous = 82;
@(negedge clk)
ifm_address_write_previous = 8'd82;
data_in_from_previous = 83;
@(negedge clk)
ifm_address_write_previous = 8'd83;
data_in_from_previous = 84;
@(negedge clk)
ifm_address_write_previous = 8'd84;
data_in_from_previous = 85;
@(negedge clk)
ifm_address_write_previous = 8'd85;
data_in_from_previous = 86;
@(negedge clk)
ifm_address_write_previous = 8'd86;
data_in_from_previous = 87;
@(negedge clk)
ifm_address_write_previous = 8'd87;
data_in_from_previous = 88;
@(negedge clk)
ifm_address_write_previous = 8'd88;
data_in_from_previous = 89;
@(negedge clk)
ifm_address_write_previous = 8'd89;
data_in_from_previous = 90;
@(negedge clk)
ifm_address_write_previous = 8'd90;
data_in_from_previous = 91;
@(negedge clk)
ifm_address_write_previous = 8'd91;
data_in_from_previous = 92;
@(negedge clk)
ifm_address_write_previous = 8'd92;
data_in_from_previous = 93;
@(negedge clk)
ifm_address_write_previous = 8'd93;
data_in_from_previous = 94;
@(negedge clk)
ifm_address_write_previous = 8'd94;
data_in_from_previous = 95;
@(negedge clk)
ifm_address_write_previous = 8'd95;
data_in_from_previous = 96;
@(negedge clk)
ifm_address_write_previous = 8'd96;
data_in_from_previous = 97;
@(negedge clk)
ifm_address_write_previous = 8'd97;
data_in_from_previous = 98;
@(negedge clk)
ifm_address_write_previous = 8'd98;
data_in_from_previous = 99;
@(negedge clk)
ifm_address_write_previous = 8'd99;
data_in_from_previous = 100;
@(negedge clk)
ifm_address_write_previous = 8'd100;
data_in_from_previous = 101;
@(negedge clk)
ifm_address_write_previous = 8'd101;
data_in_from_previous = 102;
@(negedge clk)
ifm_address_write_previous = 8'd102;
data_in_from_previous = 103;
@(negedge clk)
ifm_address_write_previous = 8'd103;
data_in_from_previous = 104;
@(negedge clk)
ifm_address_write_previous = 8'd104;
data_in_from_previous = 105;
@(negedge clk)
ifm_address_write_previous = 8'd105;
data_in_from_previous = 106;
@(negedge clk)
ifm_address_write_previous = 8'd106;
data_in_from_previous = 107;
@(negedge clk)
ifm_address_write_previous = 8'd107;
data_in_from_previous = 108;
@(negedge clk)
ifm_address_write_previous = 8'd108;
data_in_from_previous = 109;
@(negedge clk)
ifm_address_write_previous = 8'd109;
data_in_from_previous = 110;
@(negedge clk)
ifm_address_write_previous = 8'd110;
data_in_from_previous = 111;
@(negedge clk)
ifm_address_write_previous = 8'd111;
data_in_from_previous = 112;
@(negedge clk)
ifm_address_write_previous = 8'd112;
data_in_from_previous = 113;
@(negedge clk)
ifm_address_write_previous = 8'd113;
data_in_from_previous = 114;
@(negedge clk)
ifm_address_write_previous = 8'd114;
data_in_from_previous = 115;
@(negedge clk)
ifm_address_write_previous = 8'd115;
data_in_from_previous = 116;
@(negedge clk)
ifm_address_write_previous = 8'd116;
data_in_from_previous = 117;
@(negedge clk)
ifm_address_write_previous = 8'd117;
data_in_from_previous = 118;
@(negedge clk)
ifm_address_write_previous = 8'd118;
data_in_from_previous = 119;
@(negedge clk)
ifm_address_write_previous = 8'd119;
data_in_from_previous = 120;
@(negedge clk)
ifm_address_write_previous = 8'd120;
data_in_from_previous = 121;
@(negedge clk)
ifm_address_write_previous = 8'd121;
data_in_from_previous = 122;
@(negedge clk)
ifm_address_write_previous = 8'd122;
data_in_from_previous = 123;
@(negedge clk)
ifm_address_write_previous = 8'd123;
data_in_from_previous = 124;
@(negedge clk)
ifm_address_write_previous = 8'd124;
data_in_from_previous = 125;
@(negedge clk)
ifm_address_write_previous = 8'd125;
data_in_from_previous = 126;
@(negedge clk)
ifm_address_write_previous = 8'd126;
data_in_from_previous = 127;
@(negedge clk)
ifm_address_write_previous = 8'd127;
data_in_from_previous = 128;
@(negedge clk)
ifm_address_write_previous = 8'd128;
data_in_from_previous = 129;
@(negedge clk)
ifm_address_write_previous = 8'd129;
data_in_from_previous = 130;
@(negedge clk)
ifm_address_write_previous = 8'd130;
data_in_from_previous = 131;
@(negedge clk)
ifm_address_write_previous = 8'd131;
data_in_from_previous = 132;
@(negedge clk)
ifm_address_write_previous = 8'd132;
data_in_from_previous = 133;
@(negedge clk)
ifm_address_write_previous = 8'd133;
data_in_from_previous = 134;
@(negedge clk)
ifm_address_write_previous = 8'd134;
data_in_from_previous = 135;
@(negedge clk)
ifm_address_write_previous = 8'd135;
data_in_from_previous = 136;
@(negedge clk)
ifm_address_write_previous = 8'd136;
data_in_from_previous = 137;
@(negedge clk)
ifm_address_write_previous = 8'd137;
data_in_from_previous = 138;
@(negedge clk)
ifm_address_write_previous = 8'd138;
data_in_from_previous = 139;
@(negedge clk)
ifm_address_write_previous = 8'd139;
data_in_from_previous = 140;
@(negedge clk)
ifm_address_write_previous = 8'd140;
data_in_from_previous = 141;
@(negedge clk)
ifm_address_write_previous = 8'd141;
data_in_from_previous = 142;
@(negedge clk)
ifm_address_write_previous = 8'd142;
data_in_from_previous = 143;
@(negedge clk)
ifm_address_write_previous = 8'd143;
data_in_from_previous = 144;
@(negedge clk)
ifm_address_write_previous = 8'd144;
data_in_from_previous = 145;
@(negedge clk)
ifm_address_write_previous = 8'd145;
data_in_from_previous = 146;
@(negedge clk)
ifm_address_write_previous = 8'd146;
data_in_from_previous = 147;
@(negedge clk)
ifm_address_write_previous = 8'd147;
data_in_from_previous = 148;
@(negedge clk)
ifm_address_write_previous = 8'd148;
data_in_from_previous = 149;
@(negedge clk)
ifm_address_write_previous = 8'd149;
data_in_from_previous = 150;
@(negedge clk)
ifm_address_write_previous = 8'd150;
data_in_from_previous = 151;
@(negedge clk)
ifm_address_write_previous = 8'd151;
data_in_from_previous = 152;
@(negedge clk)
ifm_address_write_previous = 8'd152;
data_in_from_previous = 153;
@(negedge clk)
ifm_address_write_previous = 8'd153;
data_in_from_previous = 154;
@(negedge clk)
ifm_address_write_previous = 8'd154;
data_in_from_previous = 155;
@(negedge clk)
ifm_address_write_previous = 8'd155;
data_in_from_previous = 156;
@(negedge clk)
ifm_address_write_previous = 8'd156;
data_in_from_previous = 157;
@(negedge clk)
ifm_address_write_previous = 8'd157;
data_in_from_previous = 158;
@(negedge clk)
ifm_address_write_previous = 8'd158;
data_in_from_previous = 159;
@(negedge clk)
ifm_address_write_previous = 8'd159;
data_in_from_previous = 160;
@(negedge clk)
ifm_address_write_previous = 8'd160;
data_in_from_previous = 161;
@(negedge clk)
ifm_address_write_previous = 8'd161;
data_in_from_previous = 162;
@(negedge clk)
ifm_address_write_previous = 8'd162;
data_in_from_previous = 163;
@(negedge clk)
ifm_address_write_previous = 8'd163;
data_in_from_previous = 164;
@(negedge clk)
ifm_address_write_previous = 8'd164;
data_in_from_previous = 165;
@(negedge clk)
ifm_address_write_previous = 8'd165;
data_in_from_previous = 166;
@(negedge clk)
ifm_address_write_previous = 8'd166;
data_in_from_previous = 167;
@(negedge clk)
ifm_address_write_previous = 8'd167;
data_in_from_previous = 168;
@(negedge clk)
ifm_address_write_previous = 8'd168;
data_in_from_previous = 169;
@(negedge clk)
ifm_address_write_previous = 8'd169;
data_in_from_previous = 170;
@(negedge clk)
ifm_address_write_previous = 8'd170;
data_in_from_previous = 171;
@(negedge clk)
ifm_address_write_previous = 8'd171;
data_in_from_previous = 172;
@(negedge clk)
ifm_address_write_previous = 8'd172;
data_in_from_previous = 173;
@(negedge clk)
ifm_address_write_previous = 8'd173;
data_in_from_previous = 174;
@(negedge clk)
ifm_address_write_previous = 8'd174;
data_in_from_previous = 175;
@(negedge clk)
ifm_address_write_previous = 8'd175;
data_in_from_previous = 176;
@(negedge clk)
ifm_address_write_previous = 8'd176;
data_in_from_previous = 177;
@(negedge clk)
ifm_address_write_previous = 8'd177;
data_in_from_previous = 178;
@(negedge clk)
ifm_address_write_previous = 8'd178;
data_in_from_previous = 179;
@(negedge clk)
ifm_address_write_previous = 8'd179;
data_in_from_previous = 180;
@(negedge clk)
ifm_address_write_previous = 8'd180;
data_in_from_previous = 181;
@(negedge clk)
ifm_address_write_previous = 8'd181;
data_in_from_previous = 182;
@(negedge clk)
ifm_address_write_previous = 8'd182;
data_in_from_previous = 183;
@(negedge clk)
ifm_address_write_previous = 8'd183;
data_in_from_previous = 184;
@(negedge clk)
ifm_address_write_previous = 8'd184;
data_in_from_previous = 185;
@(negedge clk)
ifm_address_write_previous = 8'd185;
data_in_from_previous = 186;
@(negedge clk)
ifm_address_write_previous = 8'd186;
data_in_from_previous = 187;
@(negedge clk)
ifm_address_write_previous = 8'd187;
data_in_from_previous = 188;
@(negedge clk)
ifm_address_write_previous = 8'd188;
data_in_from_previous = 189;
@(negedge clk)
ifm_address_write_previous = 8'd189;
data_in_from_previous = 190;
@(negedge clk)
ifm_address_write_previous = 8'd190;
data_in_from_previous = 191;
@(negedge clk)
ifm_address_write_previous = 8'd191;
data_in_from_previous = 192;
@(negedge clk)
ifm_address_write_previous = 8'd192;
data_in_from_previous = 193;
@(negedge clk)
ifm_address_write_previous = 8'd193;
data_in_from_previous = 194;
@(negedge clk)
ifm_address_write_previous = 8'd194;
data_in_from_previous = 195;
@(negedge clk)
ifm_address_write_previous = 8'd195;
data_in_from_previous = 196;*/
/*#13900
@(negedge clk)
start_from_previous = 1'b1;
ifm_enable_write_previous = 1'b0;
@(negedge clk)
start_from_previous = 1'b0*/
end   
always #10 clk=~clk;
endmodule

